module {{cookiecutter.project_slug}} #(

)(

);
    always @() begin

    end
endmodule
